

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


package pkg is
  TYPE mem is ARRAY ( 0 to 31) of std_logic_vector( 15 downto 0);
  TYPE mem_8 is ARRAY ( 0 to 31) of std_logic_vector( 7 downto 0);
end package;

package body pkg is
end package body;
